* zero_x1
.subckt zero_x1 vdd vss zero
Mn vss one zero vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.43um
Mp one zero vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.82um
.ends zero_x1
