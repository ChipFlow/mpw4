* StdCellLib

* a2_x2
.subckt a2_x2 vss q vdd i0 i1
Mn_net0_1 vss _net0 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_net0_1 vdd _net0 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_i0_1 _net0 i0 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_i0_1 vdd i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_i1_1 _net0 i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i1_1 _net1 i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
.ends a2_x2

* a3_x2
.subckt a3_x2 vss q vdd i0 i1 i2
Mn_net1_1 vss _net1 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_net1_1 vdd _net1 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mp_i0_1 _net1 i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i0_1 _net1 i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mn_i1_1 _net0 i1 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_i1_1 vdd i1 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i2_1 _net2 i2 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_i2_1 _net1 i2 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends a3_x2

* a4_x2
.subckt a4_x2 vdd q vss i0 i1 i2 i3
Mp_net1_1 vdd _net1 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_net1_1 vss _net1 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mn_i0_1 _net1 i0 _net3 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_i0_1 vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_i1_1 _net1 i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i1_1 _net3 i1 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_i2_1 vdd i2 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i2_1 _net0 i2 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_i3_1 _net1 i3 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i3_1 _net2 i3 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
.ends a4_x2

* ao22_x2
.subckt ao22_x2 vdd q vss i0 i1 i2
Mp_net0_1 vdd _net0 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_net0_1 vss _net0 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_i0_1 vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i0_1 _net2 i0 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_i1_1 _net0 i1 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i1_1 _net1 i1 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_i2_1 _net0 i2 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i2_1 _net2 i2 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
.ends ao22_x2

* mx2_x2
.subckt mx2_x2 vdd q vss cmd i0 i1
Mp_net1_1 vdd _net1 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_net1_1 vss _net1 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_net5_1 _net1 _net5 _net4 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_net5_1 _net2 _net5 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_cmd_1 _net5 cmd vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_cmd_2 _net1 cmd _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_cmd_2 _net3 cmd _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_cmd_1 _net5 cmd vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mn_i0_1 vss i0 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_i0_1 vdd i0 _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_i1_1 _net4 i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i1_1 _net0 i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
.ends mx2_x2

* nsnrlatch_x1
.subckt nsnrlatch_x1 q vdd nq vss nrst nset
Mp_nq_1 q nq vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nq_1 _net1 nq vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_nrst_1 nq nrst vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nrst_1 _net0 nrst nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_nset_1 vdd nset q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nset_1 q nset _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp_q_1 vdd q nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_q_1 vss q _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
.ends nsnrlatch_x1

* nxr2_x1
.subckt nxr2_x1 nq vdd vss i0 i1
Mp_net0_1 nq _net0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_net0_1 nq _net0 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mn_net3_1 _net4 _net3 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_net3_1 _net1 _net3 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_i0_1 _net0 i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_i0_2 vss i0 _net4 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_i0_1 _net0 i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_i0_2 vdd i0 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mp_i1_1 _net1 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_i1_1 _net2 i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mn_i1_2 vss i1 _net3 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i1_2 vdd i1 _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends nxr2_x1

* o2_x2
.subckt o2_x2 vss q vdd i0 i1
Mn_net1_1 vss _net1 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_net1_1 vdd _net1 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mp_i0_1 _net0 i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn_i0_1 _net1 i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_i1_1 vss i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i1_1 _net1 i1 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
.ends o2_x2

* o3_x2
.subckt o3_x2 vss q vdd i0 i1 i2
Mn_net1_1 vss _net1 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_net1_1 vdd _net1 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_i0_1 _net1 i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i0_1 _net2 i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mp_i1_1 _net0 i1 _net2 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn_i1_1 vss i1 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_i2_1 _net1 i2 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i2_1 _net1 i2 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
.ends o3_x2

* o4_x2
.subckt o4_x2 vss q vdd i0 i1 i2 i3
Mn_net2_1 vss _net2 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_net2_1 vdd _net2 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_i0_1 vss i0 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i0_1 _net3 i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn_i1_1 _net2 i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i1_1 _net1 i1 _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn_i2_1 _net2 i2 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i2_1 _net0 i2 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn_i3_1 vss i3 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i3_1 _net2 i3 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
.ends o4_x2

* oa22_x2
.subckt oa22_x2 vdd q vss i0 i1 i2
Mp_net0_1 vdd _net0 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_net0_1 vss _net0 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mn_i0_1 vss i0 _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_i0_1 _net1 i0 _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i1_1 _net2 i1 _net0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_i1_1 _net0 i1 _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i2_1 _net0 i2 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_i2_1 _net1 i2 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends oa22_x2

* powmid_x0
.subckt powmid_x0 vss vdd

.ends powmid_x0

* sff1_x4
.subckt sff1_x4 vss ck vdd i q
Mn_ck nckr ck vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_ck nckr ck vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_ckr_1 _net1 ckr sff_m vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_ckr_2 y ckr sff_s vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_ckr_1 sff_m ckr _net4 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_ckr_2 sff_s ckr _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i u i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i u i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_2 sff_m nckr _net5 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_3 y nckr sff_s vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_1 vdd nckr ckr vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nckr_1 vss nckr ckr vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nckr_3 sff_s nckr _net6 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nckr_2 _net2 nckr sff_m vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_q_1 _net6 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_q_1 _net0 q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_sffm_1 vss sff_m y vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_sffm_1 vdd sff_m y vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_sffs_1 vss sff_s q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_sffs_1 vdd sff_s q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mp_sffs_2 q sff_s vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_sffs_2 q sff_s vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mn_u vss u _net2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_u vdd u _net1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_y_1 _net4 y vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_y_1 _net5 y vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends sff1_x4

* sff1r_x4
.subckt sff1r_x4 vss ck vdd i nrst q
Mn_ck_1 nckr ck vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_ck_1 nckr ck vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_ckr_1 _net0 ckr sff_m vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_ckr_2 y ckr sff_s vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_ckr_2 sff_s ckr _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_ckr_1 sff_m ckr _net6 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i_1 u i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_i_1 u i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_nckr_1 vdd nckr ckr vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nckr_1 vss nckr ckr vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nckr_2 _net7 nckr sff_m vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_nckr_3 y nckr sff_s vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nckr_2 sff_m nckr _net2 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_nckr_3 sff_s nckr _net8 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nrst_2 _net8 nrst _net5 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_nrst_1 _net4 nrst y vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_nrst_1 y nrst vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_nrst_2 vdd nrst _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_q_1 _net5 q vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_q_1 _net3 q vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_sffm_1 vdd sff_m y vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_sffm_1 vss sff_m _net4 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
Mp_sffs_1 vdd sff_s q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_sffs_2 q sff_s vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_sffs_2 q sff_s vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_sffs_1 vss sff_s q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_u_1 vdd u _net0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_u_1 vss u _net7 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_y_1 _net2 y vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn_y_1 _net6 y vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.9um
.ends sff1r_x4

* xr2_x1
.subckt xr2_x1 q vss vdd i0 i1
Mn_net0_1 q _net0 _net4 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_net0_1 q _net0 _net2 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_net3_1 _net4 _net3 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_net3_1 _net2 _net3 q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_i0_1 _net0 i0 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn_i0_2 vss i0 _net1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_i0_1 _net0 i0 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp_i0_2 vdd i0 _net2 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_i1_1 _net1 i1 q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.9um
Mp_i1_1 _net2 i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=4.0um
Mn_i1_2 vss i1 _net3 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp_i1_2 vdd i1 _net3 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends xr2_x1

* fill
.subckt fill vdd vss

.ends fill

* tie
.subckt tie vdd vss

.ends tie

* tie_diff
.subckt tie_diff vdd vss

.ends tie_diff

* tie_poly
.subckt tie_poly vdd vss

.ends tie_poly

* diode_w1
.subckt diode_w1 vdd vss i

.ends diode_w1

* zero_x1
.subckt zero_x1 vdd vss zero
Mn vss one zero vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.43um
Mp one zero vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.82um
.ends zero_x1

* one_x1
.subckt one_x1 vdd vss one
Mn vss one zero vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.43um
Mp one zero vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.82um
.ends one_x1

* zeroone_x1
.subckt zeroone_x1 vdd vss zero one
Mn vss one zero vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.43um
Mp one zero vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.82um
.ends zeroone_x1

* decap_w0
.subckt decap_w0 vdd vss
Mn vss one zero vss sky130_fd_pr__nfet_01v8__model l=0.15um w=3.43um
Mp one zero vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.82um
.ends decap_w0

* inv_x0
.subckt inv_x0 vdd vss i nq
Mn vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends inv_x0

* inv_x1
.subckt inv_x1 vdd vss i nq
Mn vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mp vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
.ends inv_x1

* inv_x2
.subckt inv_x2 vdd vss i nq
Mn0 vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mn1 nq i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mp0 vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
Mp1 nq i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
.ends inv_x2

* inv_x4
.subckt inv_x4 vdd vss i nq
Mn0 vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mn1 nq i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mn2 vss i nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mn3 nq i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mp0 vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
Mp1 nq i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
Mp2 vdd i nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
Mp3 nq i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
.ends inv_x4

* buf_x1
.subckt buf_x1 vdd vss i q
Mn1 ni i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=0.5um
Mn2_0 vss ni q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mp1 ni i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=1.0um
Mp2_0 vdd ni q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
.ends buf_x1

* buf_x2
.subckt buf_x2 vdd vss i q
Mn1 ni i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mn2_0 vss ni q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mn2_1 q ni vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mp1 ni i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mp2_0 vdd ni q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
Mp2_1 q ni vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
.ends buf_x2

* buf_x4
.subckt buf_x4 vdd vss i q
Mn1 ni i vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mn2_0 vss ni q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mn2_1 q ni vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mn2_2 vss ni q vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mn2_3 q ni vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.8um
Mp1 ni i vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
Mp2_0 vdd ni q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
Mp2_1 q ni vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
Mp2_2 vdd ni q vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
Mp2_3 q ni vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.6um
.ends buf_x4

* nand2_x0
.subckt nand2_x0 vdd vss nq i0 i1
Mn0 vss i0 int0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp0 vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
Mn1 int0 i1 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.0um
Mp1 nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.0um
.ends nand2_x0

* nand3_x0
.subckt nand3_x0 vdd vss nq i0 i1 i2
Mn0 vss i0 int0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.5um
Mp0 vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.5um
Mn1 int0 i1 int1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.5um
Mp1 nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.5um
Mn2 int1 i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.5um
Mp2 vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.5um
.ends nand3_x0

* nand4_x0
.subckt nand4_x0 vdd vss nq i0 i1 i2 i3
Mn0 vss i0 int0 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.5um
Mp0 vdd i0 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.5um
Mn1 int0 i1 int1 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.5um
Mp1 nq i1 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.5um
Mn2 int1 i2 int2 vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.5um
Mp2 vdd i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.5um
Mn3 int2 i3 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=2.5um
Mp3 nq i3 vdd vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=2.5um
.ends nand4_x0

* nor2_x0
.subckt nor2_x0 vdd vss nq i0 i1
Mn0 vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp0 vdd i0 int0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn1 nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp1 int0 i1 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
.ends nor2_x0

* nor3_x0
.subckt nor3_x0 vdd vss nq i0 i1 i2
Mn0 vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp0 vdd i0 int0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn1 nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp1 int0 i1 int1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn2 vss i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp2 int1 i2 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
.ends nor3_x0

* nor4_x0
.subckt nor4_x0 vdd vss nq i0 i1 i2 i3
Mn0 vss i0 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp0 vdd i0 int0 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn1 nq i1 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp1 int0 i1 int1 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn2 vss i2 nq vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp2 int1 i2 int2 vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
Mn3 nq i3 vss vss sky130_fd_pr__nfet_01v8__model l=0.15um w=1.0um
Mp3 int2 i3 nq vdd sky130_fd_pr__pfet_01v8__model l=0.15um w=3.0um
.ends nor4_x0
